/* 
  C6288        : Rangkaian multiplier 16x16
  Ninputs      : 32
  Noutputs     : 32
*/ 


module c6288 (
    in1,  in2,  in3,  in4,  in5,  in6,  in7,  in8, 
    in9,  in10, in11, in12, in13, in14, in15, in16,
    in17, in18, in19, in20, in21, in22, in23, in24,
    in25, in26, in27, in28, in29, in30, in31, in32,
    out1,  out2,  out3,  out4,  out5,  out6,  out7,  out8, 
    out9,  out10, out11, out12, out13, out14, out15, out16, 
    out17, out18, out19, out20, out21, out22, out23, out24, 
    out25, out26, out27, out28, out29, out30, out31, out32
);

     input  in1,  in2,  in3,  in4,  in5,  in6,  in7,  in8, 
            in9,  in10, in11, in12, in13, in14, in15, in16,
            in17, in18, in19, in20, in21, in22, in23, in24,
            in25, in26, in27, in28, in29, in30, in31, in32;

     output out1,  out2,  out3,  out4,  out5,  out6,  out7,  out8, 
            out9,  out10, out11, out12, out13, out14, out15, out16, 
            out17, out18, out19, out20, out21, out22, out23, out24, 
            out25, out26, out27, out28, out29, out30, out31, out32;

     wire [15:0] A, B;
     wire [31:0] P;

     assign
          A = {in1,  in2,  in3,  in4,  in5,  in6,  in7,  in8, 
                     in9,  in10, in11, in12, in13, in14, in15, in16},
      
          B = {in17, in18, in19, in20, in21, in22, in23, in24,
                     in25, in26, in27, in28, in29, in30, in31, in32},

          {out1,  out2,  out3,  out4,  out5,  out6,  out7,  out8, 
          out9,  out10, out11, out12, out13, out14, out15, out16, 
          out17, out18, out19, out20, out21, out22, out23, out24, 
          out25, out26, out27, out28, out29, out30, out31, out32} 
          = P;

     assign P = A * B;
endmodule 